** sch_path: /home/hoyeon/Desktop/ciropt/netlist/simplecsamp
**.subckt simplecsamp
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L = {Length1}  W = {Width1} nf = {Nf1} ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V3 net1 GND 0
V4 net2 GND 0.9
**** begin user architecture code
** design_variables_start
.param Length1 = 0.15
.param Width1 = 1
.param Nf1 = 1

** design_variables_end
.lib /home/hoyeon/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.control
	dc V3 0 3 0.01
.endc

.save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
